-- megafunction wizard: %Arria V Transceiver Native PHY v15.1%
-- GENERATION: XML
-- GXB_RX.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity GXB_RX is
	port (
		rx_analogreset          : in  std_logic_vector(3 downto 0)   := (others => '0'); --          rx_analogreset.rx_analogreset
		rx_digitalreset         : in  std_logic_vector(3 downto 0)   := (others => '0'); --         rx_digitalreset.rx_digitalreset
		rx_cdr_refclk           : in  std_logic_vector(0 downto 0)   := (others => '0'); --           rx_cdr_refclk.rx_cdr_refclk
		rx_serial_data          : in  std_logic_vector(3 downto 0)   := (others => '0'); --          rx_serial_data.rx_serial_data
		rx_std_coreclkin        : in  std_logic_vector(3 downto 0)   := (others => '0'); --        rx_std_coreclkin.rx_std_coreclkin
		rx_std_clkout           : out std_logic_vector(3 downto 0);                      --           rx_std_clkout.rx_std_clkout
		rx_cal_busy             : out std_logic_vector(3 downto 0);                      --             rx_cal_busy.rx_cal_busy
		reconfig_to_xcvr        : in  std_logic_vector(279 downto 0) := (others => '0'); --        reconfig_to_xcvr.reconfig_to_xcvr
		reconfig_from_xcvr      : out std_logic_vector(183 downto 0);                    --      reconfig_from_xcvr.reconfig_from_xcvr
		rx_parallel_data        : out std_logic_vector(63 downto 0);                     --        rx_parallel_data.rx_parallel_data
		rx_datak                : out std_logic_vector(7 downto 0);                      --                rx_datak.rx_datak
		rx_errdetect            : out std_logic_vector(7 downto 0);                      --            rx_errdetect.rx_errdetect
		rx_disperr              : out std_logic_vector(7 downto 0);                      --              rx_disperr.rx_disperr
		rx_runningdisp          : out std_logic_vector(7 downto 0);                      --          rx_runningdisp.rx_runningdisp
		rx_patterndetect        : out std_logic_vector(7 downto 0);                      --        rx_patterndetect.rx_patterndetect
		rx_syncstatus           : out std_logic_vector(7 downto 0);                      --           rx_syncstatus.rx_syncstatus
		unused_rx_parallel_data : out std_logic_vector(143 downto 0)                     -- unused_rx_parallel_data.unused_rx_parallel_data
	);
end entity GXB_RX;

architecture rtl of GXB_RX is
	component altera_xcvr_native_av is
		generic (
			tx_enable                       : integer := 1;
			rx_enable                       : integer := 1;
			enable_std                      : integer := 0;
			data_path_select                : string  := "pma_direct";
			channels                        : integer := 1;
			bonded_mode                     : string  := "non_bonded";
			data_rate                       : string  := "";
			pma_width                       : integer := 80;
			tx_pma_clk_div                  : integer := 1;
			pll_reconfig_enable             : integer := 0;
			pll_external_enable             : integer := 0;
			pll_data_rate                   : string  := "0 Mbps";
			pll_type                        : string  := "CMU";
			pma_bonding_mode                : string  := "x1";
			plls                            : integer := 1;
			pll_select                      : integer := 0;
			pll_refclk_cnt                  : integer := 1;
			pll_refclk_select               : string  := "0";
			pll_refclk_freq                 : string  := "125.0 MHz";
			pll_feedback_path               : string  := "internal";
			cdr_reconfig_enable             : integer := 0;
			cdr_refclk_cnt                  : integer := 1;
			cdr_refclk_select               : integer := 0;
			cdr_refclk_freq                 : string  := "";
			rx_ppm_detect_threshold         : string  := "1000";
			rx_clkslip_enable               : integer := 0;
			std_protocol_hint               : string  := "basic";
			std_pcs_pma_width               : integer := 10;
			std_low_latency_bypass_enable   : integer := 0;
			std_tx_pcfifo_mode              : string  := "low_latency";
			std_rx_pcfifo_mode              : string  := "low_latency";
			std_rx_byte_order_enable        : integer := 0;
			std_rx_byte_order_mode          : string  := "manual";
			std_rx_byte_order_width         : integer := 10;
			std_rx_byte_order_symbol_count  : integer := 1;
			std_rx_byte_order_pattern       : string  := "0";
			std_rx_byte_order_pad           : string  := "0";
			std_tx_byte_ser_enable          : integer := 0;
			std_rx_byte_deser_enable        : integer := 0;
			std_tx_8b10b_enable             : integer := 0;
			std_tx_8b10b_disp_ctrl_enable   : integer := 0;
			std_rx_8b10b_enable             : integer := 0;
			std_rx_rmfifo_enable            : integer := 0;
			std_rx_rmfifo_pattern_p         : string  := "00000";
			std_rx_rmfifo_pattern_n         : string  := "00000";
			std_tx_bitslip_enable           : integer := 0;
			std_rx_word_aligner_mode        : string  := "bit_slip";
			std_rx_word_aligner_pattern_len : integer := 7;
			std_rx_word_aligner_pattern     : string  := "0000000000";
			std_rx_word_aligner_rknumber    : integer := 3;
			std_rx_word_aligner_renumber    : integer := 3;
			std_rx_word_aligner_rgnumber    : integer := 3;
			std_rx_run_length_val           : integer := 31;
			std_tx_bitrev_enable            : integer := 0;
			std_rx_bitrev_enable            : integer := 0;
			std_tx_byterev_enable           : integer := 0;
			std_rx_byterev_enable           : integer := 0;
			std_tx_polinv_enable            : integer := 0;
			std_rx_polinv_enable            : integer := 0
		);
		port (
			rx_analogreset            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_digitalreset
			rx_cdr_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- rx_cdr_refclk
			rx_serial_data            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_std_coreclkin          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_coreclkin
			rx_std_clkout             : out std_logic_vector(3 downto 0);                      -- rx_std_clkout
			rx_cal_busy               : out std_logic_vector(3 downto 0);                      -- rx_cal_busy
			reconfig_to_xcvr          : in  std_logic_vector(279 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			reconfig_from_xcvr        : out std_logic_vector(183 downto 0);                    -- reconfig_from_xcvr
			rx_parallel_data          : out std_logic_vector(255 downto 0);                    -- unused_rx_parallel_data
			pll_powerdown             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- pll_powerdown
			tx_analogreset            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_digitalreset
			tx_pll_refclk             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_pll_refclk
			tx_pma_clkout             : out std_logic_vector(3 downto 0);                      -- tx_pma_clkout
			tx_serial_data            : out std_logic_vector(3 downto 0);                      -- tx_serial_data
			tx_pma_parallel_data      : in  std_logic_vector(319 downto 0) := (others => 'X'); -- tx_pma_parallel_data
			pll_locked                : out std_logic_vector(3 downto 0);                      -- pll_locked
			ext_pll_clk               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- ext_pll_clk
			rx_pma_clkout             : out std_logic_vector(3 downto 0);                      -- rx_pma_clkout
			rx_pma_parallel_data      : out std_logic_vector(319 downto 0);                    -- rx_pma_parallel_data
			rx_clkslip                : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_clkslip
			rx_clklow                 : out std_logic_vector(3 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(3 downto 0);                      -- rx_fref
			rx_set_locktodata         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_is_lockedtoref         : out std_logic_vector(3 downto 0);                      -- rx_is_lockedtoref
			rx_is_lockedtodata        : out std_logic_vector(3 downto 0);                      -- rx_is_lockedtodata
			rx_seriallpbken           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_seriallpbken
			rx_signaldetect           : out std_logic_vector(3 downto 0);                      -- rx_signaldetect
			tx_parallel_data          : in  std_logic_vector(175 downto 0) := (others => 'X'); -- tx_parallel_data
			tx_std_coreclkin          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_std_coreclkin
			tx_std_clkout             : out std_logic_vector(3 downto 0);                      -- tx_std_clkout
			rx_std_prbs_done          : out std_logic_vector(3 downto 0);                      -- rx_std_prbs_done
			rx_std_prbs_err           : out std_logic_vector(3 downto 0);                      -- rx_std_prbs_err
			tx_std_pcfifo_full        : out std_logic_vector(3 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(3 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(3 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(3 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_byteorder_ena      : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_byteorder_ena
			rx_std_byteorder_flag     : out std_logic_vector(3 downto 0);                      -- rx_std_byteorder_flag
			rx_std_rmfifo_full        : out std_logic_vector(3 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(3 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_wa_patternalign    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			rx_std_wa_a1a2size        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			tx_std_bitslipboundarysel : in  std_logic_vector(19 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(19 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_bitslip            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_bitslip
			rx_std_runlength_err      : out std_logic_vector(3 downto 0);                      -- rx_std_runlength_err
			rx_std_bitrev_ena         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_std_polinv             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_std_polinv
			rx_std_polinv             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_polinv
			tx_std_elecidle           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_std_elecidle
			rx_std_signaldetect       : out std_logic_vector(3 downto 0);                      -- rx_std_signaldetect
			tx_cal_busy               : out std_logic_vector(3 downto 0)                       -- tx_cal_busy
		);
	end component altera_xcvr_native_av;

	signal gxb_rx_inst_rx_parallel_data : std_logic_vector(255 downto 0); -- port fragment

begin

	gxb_rx_inst : component altera_xcvr_native_av
		generic map (
			tx_enable                       => 0,
			rx_enable                       => 1,
			enable_std                      => 1,
			data_path_select                => "standard",
			channels                        => 4,
			bonded_mode                     => "non_bonded",
			data_rate                       => "1280 Mbps",
			pma_width                       => 10,
			tx_pma_clk_div                  => 1,
			pll_reconfig_enable             => 0,
			pll_external_enable             => 0,
			pll_data_rate                   => "1280 Mbps",
			pll_type                        => "CMU",
			pma_bonding_mode                => "x1",
			plls                            => 1,
			pll_select                      => 0,
			pll_refclk_cnt                  => 1,
			pll_refclk_select               => "0",
			pll_refclk_freq                 => "unused",
			pll_feedback_path               => "internal",
			cdr_reconfig_enable             => 0,
			cdr_refclk_cnt                  => 1,
			cdr_refclk_select               => 0,
			cdr_refclk_freq                 => "128.0 MHz",
			rx_ppm_detect_threshold         => "1000",
			rx_clkslip_enable               => 0,
			std_protocol_hint               => "basic",
			std_pcs_pma_width               => 10,
			std_low_latency_bypass_enable   => 0,
			std_tx_pcfifo_mode              => "low_latency",
			std_rx_pcfifo_mode              => "register_fifo",
			std_rx_byte_order_enable        => 1,
			std_rx_byte_order_mode          => "auto",
			std_rx_byte_order_width         => 9,
			std_rx_byte_order_symbol_count  => 1,
			std_rx_byte_order_pattern       => "1fb",
			std_rx_byte_order_pad           => "0",
			std_tx_byte_ser_enable          => 0,
			std_rx_byte_deser_enable        => 1,
			std_tx_8b10b_enable             => 0,
			std_tx_8b10b_disp_ctrl_enable   => 0,
			std_rx_8b10b_enable             => 1,
			std_rx_rmfifo_enable            => 0,
			std_rx_rmfifo_pattern_p         => "00000",
			std_rx_rmfifo_pattern_n         => "00000",
			std_tx_bitslip_enable           => 0,
			std_rx_word_aligner_mode        => "sync_sm",
			std_rx_word_aligner_pattern_len => 10,
			std_rx_word_aligner_pattern     => "17c",
			std_rx_word_aligner_rknumber    => 2,
			std_rx_word_aligner_renumber    => 3,
			std_rx_word_aligner_rgnumber    => 3,
			std_rx_run_length_val           => 2,
			std_tx_bitrev_enable            => 0,
			std_rx_bitrev_enable            => 0,
			std_tx_byterev_enable           => 0,
			std_rx_byterev_enable           => 0,
			std_tx_polinv_enable            => 0,
			std_rx_polinv_enable            => 0
		)
		port map (
			rx_analogreset            => rx_analogreset,                                                                                                                                                                                                                                                                                                                     --     rx_analogreset.rx_analogreset
			rx_digitalreset           => rx_digitalreset,                                                                                                                                                                                                                                                                                                                    --    rx_digitalreset.rx_digitalreset
			rx_cdr_refclk             => rx_cdr_refclk,                                                                                                                                                                                                                                                                                                                      --      rx_cdr_refclk.rx_cdr_refclk
			rx_serial_data            => rx_serial_data,                                                                                                                                                                                                                                                                                                                     --     rx_serial_data.rx_serial_data
			rx_std_coreclkin          => rx_std_coreclkin,                                                                                                                                                                                                                                                                                                                   --   rx_std_coreclkin.rx_std_coreclkin
			rx_std_clkout             => rx_std_clkout,                                                                                                                                                                                                                                                                                                                      --      rx_std_clkout.rx_std_clkout
			rx_cal_busy               => rx_cal_busy,                                                                                                                                                                                                                                                                                                                        --        rx_cal_busy.rx_cal_busy
			reconfig_to_xcvr          => reconfig_to_xcvr,                                                                                                                                                                                                                                                                                                                   --   reconfig_to_xcvr.reconfig_to_xcvr
			reconfig_from_xcvr        => reconfig_from_xcvr,                                                                                                                                                                                                                                                                                                                 -- reconfig_from_xcvr.reconfig_from_xcvr
			rx_parallel_data          => gxb_rx_inst_rx_parallel_data,                                                                                                                                                                                                                                                                                                       --   rx_parallel_data.rx_parallel_data
			pll_powerdown             => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_analogreset            => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_digitalreset           => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_pll_refclk             => "0",                                                                                                                                                                                                                                                                                                                                --        (terminated)
			tx_pma_clkout             => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_serial_data            => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_pma_parallel_data      => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --        (terminated)
			pll_locked                => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			ext_pll_clk               => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_pma_clkout             => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_pma_parallel_data      => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_clkslip                => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_clklow                 => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_fref                   => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_set_locktodata         => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_set_locktoref          => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_is_lockedtoref         => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_is_lockedtodata        => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_seriallpbken           => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_signaldetect           => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_parallel_data          => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",                                                                                                                                                 --        (terminated)
			tx_std_coreclkin          => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_std_clkout             => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_done          => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_prbs_err           => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_byteorder_ena      => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_byteorder_flag     => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_full        => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_rmfifo_empty       => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_wa_patternalign    => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_wa_a1a2size        => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_std_bitslipboundarysel => "00000000000000000000",                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_bitslipboundarysel => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitslip            => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_runlength_err      => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			rx_std_bitrev_ena         => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_byterev_ena        => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_std_polinv             => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_polinv             => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			tx_std_elecidle           => "0000",                                                                                                                                                                                                                                                                                                                             --        (terminated)
			rx_std_signaldetect       => open,                                                                                                                                                                                                                                                                                                                               --        (terminated)
			tx_cal_busy               => open                                                                                                                                                                                                                                                                                                                                --        (terminated)
		);

	rx_datak <= GXB_RX_inst_rx_parallel_data(232 downto 232) & GXB_RX_inst_rx_parallel_data(200 downto 200) & GXB_RX_inst_rx_parallel_data(168 downto 168) & GXB_RX_inst_rx_parallel_data(136 downto 136) & GXB_RX_inst_rx_parallel_data(104 downto 104) & GXB_RX_inst_rx_parallel_data(72 downto 72) & GXB_RX_inst_rx_parallel_data(40 downto 40) & GXB_RX_inst_rx_parallel_data(8 downto 8);

	unused_rx_parallel_data <= GXB_RX_inst_rx_parallel_data(255 downto 255) & GXB_RX_inst_rx_parallel_data(254 downto 254) & GXB_RX_inst_rx_parallel_data(253 downto 253) & GXB_RX_inst_rx_parallel_data(252 downto 252) & GXB_RX_inst_rx_parallel_data(251 downto 251) & GXB_RX_inst_rx_parallel_data(250 downto 250) & GXB_RX_inst_rx_parallel_data(249 downto 249) & GXB_RX_inst_rx_parallel_data(248 downto 248) & GXB_RX_inst_rx_parallel_data(247 downto 247) & GXB_RX_inst_rx_parallel_data(246 downto 246) & GXB_RX_inst_rx_parallel_data(245 downto 245) & GXB_RX_inst_rx_parallel_data(244 downto 244) & GXB_RX_inst_rx_parallel_data(243 downto 243) & GXB_RX_inst_rx_parallel_data(242 downto 242) & GXB_RX_inst_rx_parallel_data(241 downto 241) & GXB_RX_inst_rx_parallel_data(240 downto 240) & GXB_RX_inst_rx_parallel_data(238 downto 238) & GXB_RX_inst_rx_parallel_data(237 downto 237) & GXB_RX_inst_rx_parallel_data(223 downto 223) & GXB_RX_inst_rx_parallel_data(222 downto 222) & GXB_RX_inst_rx_parallel_data(221 downto 221) & GXB_RX_inst_rx_parallel_data(220 downto 220) & GXB_RX_inst_rx_parallel_data(219 downto 219) & GXB_RX_inst_rx_parallel_data(218 downto 218) & GXB_RX_inst_rx_parallel_data(217 downto 217) & GXB_RX_inst_rx_parallel_data(216 downto 216) & GXB_RX_inst_rx_parallel_data(215 downto 215) & GXB_RX_inst_rx_parallel_data(214 downto 214) & GXB_RX_inst_rx_parallel_data(213 downto 213) & GXB_RX_inst_rx_parallel_data(212 downto 212) & GXB_RX_inst_rx_parallel_data(211 downto 211) & GXB_RX_inst_rx_parallel_data(210 downto 210) & GXB_RX_inst_rx_parallel_data(209 downto 209) & GXB_RX_inst_rx_parallel_data(208 downto 208) & GXB_RX_inst_rx_parallel_data(206 downto 206) & GXB_RX_inst_rx_parallel_data(205 downto 205) & GXB_RX_inst_rx_parallel_data(191 downto 191) & GXB_RX_inst_rx_parallel_data(190 downto 190) & GXB_RX_inst_rx_parallel_data(189 downto 189) & GXB_RX_inst_rx_parallel_data(188 downto 188) & GXB_RX_inst_rx_parallel_data(187 downto 187) & GXB_RX_inst_rx_parallel_data(186 downto 186) & GXB_RX_inst_rx_parallel_data(185 downto 185) & GXB_RX_inst_rx_parallel_data(184 downto 184) & GXB_RX_inst_rx_parallel_data(183 downto 183) & GXB_RX_inst_rx_parallel_data(182 downto 182) & GXB_RX_inst_rx_parallel_data(181 downto 181) & GXB_RX_inst_rx_parallel_data(180 downto 180) & GXB_RX_inst_rx_parallel_data(179 downto 179) & GXB_RX_inst_rx_parallel_data(178 downto 178) & GXB_RX_inst_rx_parallel_data(177 downto 177) & GXB_RX_inst_rx_parallel_data(176 downto 176) & GXB_RX_inst_rx_parallel_data(174 downto 174) & GXB_RX_inst_rx_parallel_data(173 downto 173) & GXB_RX_inst_rx_parallel_data(159 downto 159) & GXB_RX_inst_rx_parallel_data(158 downto 158) & GXB_RX_inst_rx_parallel_data(157 downto 157) & GXB_RX_inst_rx_parallel_data(156 downto 156) & GXB_RX_inst_rx_parallel_data(155 downto 155) & GXB_RX_inst_rx_parallel_data(154 downto 154) & GXB_RX_inst_rx_parallel_data(153 downto 153) & GXB_RX_inst_rx_parallel_data(152 downto 152) & GXB_RX_inst_rx_parallel_data(151 downto 151) & GXB_RX_inst_rx_parallel_data(150 downto 150) & GXB_RX_inst_rx_parallel_data(149 downto 149) & GXB_RX_inst_rx_parallel_data(148 downto 148) & GXB_RX_inst_rx_parallel_data(147 downto 147) & GXB_RX_inst_rx_parallel_data(146 downto 146) & GXB_RX_inst_rx_parallel_data(145 downto 145) & GXB_RX_inst_rx_parallel_data(144 downto 144) & GXB_RX_inst_rx_parallel_data(142 downto 142) & GXB_RX_inst_rx_parallel_data(141 downto 141) & GXB_RX_inst_rx_parallel_data(127 downto 127) & GXB_RX_inst_rx_parallel_data(126 downto 126) & GXB_RX_inst_rx_parallel_data(125 downto 125) & GXB_RX_inst_rx_parallel_data(124 downto 124) & GXB_RX_inst_rx_parallel_data(123 downto 123) & GXB_RX_inst_rx_parallel_data(122 downto 122) & GXB_RX_inst_rx_parallel_data(121 downto 121) & GXB_RX_inst_rx_parallel_data(120 downto 120) & GXB_RX_inst_rx_parallel_data(119 downto 119) & GXB_RX_inst_rx_parallel_data(118 downto 118) & GXB_RX_inst_rx_parallel_data(117 downto 117) & GXB_RX_inst_rx_parallel_data(116 downto 116) & GXB_RX_inst_rx_parallel_data(115 downto 115) & GXB_RX_inst_rx_parallel_data(114 downto 114) & GXB_RX_inst_rx_parallel_data(113 downto 113) & GXB_RX_inst_rx_parallel_data(112 downto 112) & GXB_RX_inst_rx_parallel_data(110 downto 110) & GXB_RX_inst_rx_parallel_data(109 downto 109) & GXB_RX_inst_rx_parallel_data(95 downto 95) & GXB_RX_inst_rx_parallel_data(94 downto 94) & GXB_RX_inst_rx_parallel_data(93 downto 93) & GXB_RX_inst_rx_parallel_data(92 downto 92) & GXB_RX_inst_rx_parallel_data(91 downto 91) & GXB_RX_inst_rx_parallel_data(90 downto 90) & GXB_RX_inst_rx_parallel_data(89 downto 89) & GXB_RX_inst_rx_parallel_data(88 downto 88) & GXB_RX_inst_rx_parallel_data(87 downto 87) & GXB_RX_inst_rx_parallel_data(86 downto 86) & GXB_RX_inst_rx_parallel_data(85 downto 85) & GXB_RX_inst_rx_parallel_data(84 downto 84) & GXB_RX_inst_rx_parallel_data(83 downto 83) & GXB_RX_inst_rx_parallel_data(82 downto 82) & GXB_RX_inst_rx_parallel_data(81 downto 81) & GXB_RX_inst_rx_parallel_data(80 downto 80) & GXB_RX_inst_rx_parallel_data(78 downto 78) & GXB_RX_inst_rx_parallel_data(77 downto 77) & GXB_RX_inst_rx_parallel_data(63 downto 63) & GXB_RX_inst_rx_parallel_data(62 downto 62) & GXB_RX_inst_rx_parallel_data(61 downto 61) & GXB_RX_inst_rx_parallel_data(60 downto 60) & GXB_RX_inst_rx_parallel_data(59 downto 59) & GXB_RX_inst_rx_parallel_data(58 downto 58) & GXB_RX_inst_rx_parallel_data(57 downto 57) & GXB_RX_inst_rx_parallel_data(56 downto 56) & GXB_RX_inst_rx_parallel_data(55 downto 55) & GXB_RX_inst_rx_parallel_data(54 downto 54) & GXB_RX_inst_rx_parallel_data(53 downto 53) & GXB_RX_inst_rx_parallel_data(52 downto 52) & GXB_RX_inst_rx_parallel_data(51 downto 51) & GXB_RX_inst_rx_parallel_data(50 downto 50) & GXB_RX_inst_rx_parallel_data(49 downto 49) & GXB_RX_inst_rx_parallel_data(48 downto 48) & GXB_RX_inst_rx_parallel_data(46 downto 46) & GXB_RX_inst_rx_parallel_data(45 downto 45) & GXB_RX_inst_rx_parallel_data(31 downto 31) & GXB_RX_inst_rx_parallel_data(30 downto 30) & GXB_RX_inst_rx_parallel_data(29 downto 29) & GXB_RX_inst_rx_parallel_data(28 downto 28) & GXB_RX_inst_rx_parallel_data(27 downto 27) & GXB_RX_inst_rx_parallel_data(26 downto 26) & GXB_RX_inst_rx_parallel_data(25 downto 25) & GXB_RX_inst_rx_parallel_data(24 downto 24) & GXB_RX_inst_rx_parallel_data(23 downto 23) & GXB_RX_inst_rx_parallel_data(22 downto 22) & GXB_RX_inst_rx_parallel_data(21 downto 21) & GXB_RX_inst_rx_parallel_data(20 downto 20) & GXB_RX_inst_rx_parallel_data(19 downto 19) & GXB_RX_inst_rx_parallel_data(18 downto 18) & GXB_RX_inst_rx_parallel_data(17 downto 17) & GXB_RX_inst_rx_parallel_data(16 downto 16) & GXB_RX_inst_rx_parallel_data(14 downto 14) & GXB_RX_inst_rx_parallel_data(13 downto 13);

	rx_syncstatus <= GXB_RX_inst_rx_parallel_data(234 downto 234) & GXB_RX_inst_rx_parallel_data(202 downto 202) & GXB_RX_inst_rx_parallel_data(170 downto 170) & GXB_RX_inst_rx_parallel_data(138 downto 138) & GXB_RX_inst_rx_parallel_data(106 downto 106) & GXB_RX_inst_rx_parallel_data(74 downto 74) & GXB_RX_inst_rx_parallel_data(42 downto 42) & GXB_RX_inst_rx_parallel_data(10 downto 10);

	rx_patterndetect <= GXB_RX_inst_rx_parallel_data(236 downto 236) & GXB_RX_inst_rx_parallel_data(204 downto 204) & GXB_RX_inst_rx_parallel_data(172 downto 172) & GXB_RX_inst_rx_parallel_data(140 downto 140) & GXB_RX_inst_rx_parallel_data(108 downto 108) & GXB_RX_inst_rx_parallel_data(76 downto 76) & GXB_RX_inst_rx_parallel_data(44 downto 44) & GXB_RX_inst_rx_parallel_data(12 downto 12);

	rx_runningdisp <= GXB_RX_inst_rx_parallel_data(239 downto 239) & GXB_RX_inst_rx_parallel_data(207 downto 207) & GXB_RX_inst_rx_parallel_data(175 downto 175) & GXB_RX_inst_rx_parallel_data(143 downto 143) & GXB_RX_inst_rx_parallel_data(111 downto 111) & GXB_RX_inst_rx_parallel_data(79 downto 79) & GXB_RX_inst_rx_parallel_data(47 downto 47) & GXB_RX_inst_rx_parallel_data(15 downto 15);

	rx_parallel_data <= GXB_RX_inst_rx_parallel_data(231 downto 231) & GXB_RX_inst_rx_parallel_data(230 downto 230) & GXB_RX_inst_rx_parallel_data(229 downto 229) & GXB_RX_inst_rx_parallel_data(228 downto 228) & GXB_RX_inst_rx_parallel_data(227 downto 227) & GXB_RX_inst_rx_parallel_data(226 downto 226) & GXB_RX_inst_rx_parallel_data(225 downto 225) & GXB_RX_inst_rx_parallel_data(224 downto 224) & GXB_RX_inst_rx_parallel_data(199 downto 199) & GXB_RX_inst_rx_parallel_data(198 downto 198) & GXB_RX_inst_rx_parallel_data(197 downto 197) & GXB_RX_inst_rx_parallel_data(196 downto 196) & GXB_RX_inst_rx_parallel_data(195 downto 195) & GXB_RX_inst_rx_parallel_data(194 downto 194) & GXB_RX_inst_rx_parallel_data(193 downto 193) & GXB_RX_inst_rx_parallel_data(192 downto 192) & GXB_RX_inst_rx_parallel_data(167 downto 167) & GXB_RX_inst_rx_parallel_data(166 downto 166) & GXB_RX_inst_rx_parallel_data(165 downto 165) & GXB_RX_inst_rx_parallel_data(164 downto 164) & GXB_RX_inst_rx_parallel_data(163 downto 163) & GXB_RX_inst_rx_parallel_data(162 downto 162) & GXB_RX_inst_rx_parallel_data(161 downto 161) & GXB_RX_inst_rx_parallel_data(160 downto 160) & GXB_RX_inst_rx_parallel_data(135 downto 135) & GXB_RX_inst_rx_parallel_data(134 downto 134) & GXB_RX_inst_rx_parallel_data(133 downto 133) & GXB_RX_inst_rx_parallel_data(132 downto 132) & GXB_RX_inst_rx_parallel_data(131 downto 131) & GXB_RX_inst_rx_parallel_data(130 downto 130) & GXB_RX_inst_rx_parallel_data(129 downto 129) & GXB_RX_inst_rx_parallel_data(128 downto 128) & GXB_RX_inst_rx_parallel_data(103 downto 103) & GXB_RX_inst_rx_parallel_data(102 downto 102) & GXB_RX_inst_rx_parallel_data(101 downto 101) & GXB_RX_inst_rx_parallel_data(100 downto 100) & GXB_RX_inst_rx_parallel_data(99 downto 99) & GXB_RX_inst_rx_parallel_data(98 downto 98) & GXB_RX_inst_rx_parallel_data(97 downto 97) & GXB_RX_inst_rx_parallel_data(96 downto 96) & GXB_RX_inst_rx_parallel_data(71 downto 71) & GXB_RX_inst_rx_parallel_data(70 downto 70) & GXB_RX_inst_rx_parallel_data(69 downto 69) & GXB_RX_inst_rx_parallel_data(68 downto 68) & GXB_RX_inst_rx_parallel_data(67 downto 67) & GXB_RX_inst_rx_parallel_data(66 downto 66) & GXB_RX_inst_rx_parallel_data(65 downto 65) & GXB_RX_inst_rx_parallel_data(64 downto 64) & GXB_RX_inst_rx_parallel_data(39 downto 39) & GXB_RX_inst_rx_parallel_data(38 downto 38) & GXB_RX_inst_rx_parallel_data(37 downto 37) & GXB_RX_inst_rx_parallel_data(36 downto 36) & GXB_RX_inst_rx_parallel_data(35 downto 35) & GXB_RX_inst_rx_parallel_data(34 downto 34) & GXB_RX_inst_rx_parallel_data(33 downto 33) & GXB_RX_inst_rx_parallel_data(32 downto 32) & GXB_RX_inst_rx_parallel_data(7 downto 7) & GXB_RX_inst_rx_parallel_data(6 downto 6) & GXB_RX_inst_rx_parallel_data(5 downto 5) & GXB_RX_inst_rx_parallel_data(4 downto 4) & GXB_RX_inst_rx_parallel_data(3 downto 3) & GXB_RX_inst_rx_parallel_data(2 downto 2) & GXB_RX_inst_rx_parallel_data(1 downto 1) & GXB_RX_inst_rx_parallel_data(0 downto 0);

	rx_errdetect <= GXB_RX_inst_rx_parallel_data(233 downto 233) & GXB_RX_inst_rx_parallel_data(201 downto 201) & GXB_RX_inst_rx_parallel_data(169 downto 169) & GXB_RX_inst_rx_parallel_data(137 downto 137) & GXB_RX_inst_rx_parallel_data(105 downto 105) & GXB_RX_inst_rx_parallel_data(73 downto 73) & GXB_RX_inst_rx_parallel_data(41 downto 41) & GXB_RX_inst_rx_parallel_data(9 downto 9);

	rx_disperr <= GXB_RX_inst_rx_parallel_data(235 downto 235) & GXB_RX_inst_rx_parallel_data(203 downto 203) & GXB_RX_inst_rx_parallel_data(171 downto 171) & GXB_RX_inst_rx_parallel_data(139 downto 139) & GXB_RX_inst_rx_parallel_data(107 downto 107) & GXB_RX_inst_rx_parallel_data(75 downto 75) & GXB_RX_inst_rx_parallel_data(43 downto 43) & GXB_RX_inst_rx_parallel_data(11 downto 11);

end architecture rtl; -- of GXB_RX
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_xcvr_native_av" version="15.1" >
-- Retrieval info: 	<generic name="device_family" value="Arria V" />
-- Retrieval info: 	<generic name="show_advanced_features" value="0" />
-- Retrieval info: 	<generic name="device_speedgrade" value="fastest" />
-- Retrieval info: 	<generic name="message_level" value="error" />
-- Retrieval info: 	<generic name="tx_enable" value="0" />
-- Retrieval info: 	<generic name="rx_enable" value="1" />
-- Retrieval info: 	<generic name="enable_std" value="1" />
-- Retrieval info: 	<generic name="set_data_path_select" value="standard" />
-- Retrieval info: 	<generic name="channels" value="4" />
-- Retrieval info: 	<generic name="bonded_mode" value="non_bonded" />
-- Retrieval info: 	<generic name="enable_simple_interface" value="1" />
-- Retrieval info: 	<generic name="set_data_rate" value="1280" />
-- Retrieval info: 	<generic name="pma_direct_width" value="80" />
-- Retrieval info: 	<generic name="tx_pma_clk_div" value="1" />
-- Retrieval info: 	<generic name="pll_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="pll_external_enable" value="0" />
-- Retrieval info: 	<generic name="plls" value="1" />
-- Retrieval info: 	<generic name="pll_select" value="0" />
-- Retrieval info: 	<generic name="pll_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_reconfig_enable" value="0" />
-- Retrieval info: 	<generic name="cdr_refclk_cnt" value="1" />
-- Retrieval info: 	<generic name="cdr_refclk_select" value="0" />
-- Retrieval info: 	<generic name="set_cdr_refclk_freq" value="128.0 MHz" />
-- Retrieval info: 	<generic name="rx_ppm_detect_threshold" value="1000" />
-- Retrieval info: 	<generic name="enable_port_rx_pma_clkout" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtodata" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_is_lockedtoref" value="0" />
-- Retrieval info: 	<generic name="enable_ports_rx_manual_cdr_mode" value="0" />
-- Retrieval info: 	<generic name="rx_clkslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_seriallpbken" value="0" />
-- Retrieval info: 	<generic name="std_protocol_hint" value="basic" />
-- Retrieval info: 	<generic name="std_pcs_pma_width" value="10" />
-- Retrieval info: 	<generic name="std_low_latency_bypass_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_pcfifo_mode" value="low_latency" />
-- Retrieval info: 	<generic name="std_rx_pcfifo_mode" value="register_fifo" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_order_enable" value="1" />
-- Retrieval info: 	<generic name="std_rx_byte_order_mode" value="auto" />
-- Retrieval info: 	<generic name="std_rx_byte_order_symbol_count" value="1" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pattern" value="1fb" />
-- Retrieval info: 	<generic name="std_rx_byte_order_pad" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byteorder_flag" value="0" />
-- Retrieval info: 	<generic name="std_tx_byte_ser_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byte_deser_enable" value="1" />
-- Retrieval info: 	<generic name="std_tx_8b10b_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_8b10b_disp_ctrl_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_8b10b_enable" value="1" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_p" value="00000" />
-- Retrieval info: 	<generic name="std_rx_rmfifo_pattern_n" value="00000" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_full" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_empty" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitslip_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_mode" value="sync_sm" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern_len" value="10" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_pattern" value="17c" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rknumber" value="2" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_renumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_word_aligner_rgnumber" value="3" />
-- Retrieval info: 	<generic name="std_rx_run_length_val" value="2" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_patternalign" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_wa_a1a2size" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslipboundarysel" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitslip" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_runlength_err" value="0" />
-- Retrieval info: 	<generic name="std_tx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_bitrev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_byterev_enable" value="0" />
-- Retrieval info: 	<generic name="std_tx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="std_rx_polinv_enable" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_bitrev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_byterev_ena" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_polinv" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_polinv" value="0" />
-- Retrieval info: 	<generic name="enable_port_tx_std_elecidle" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_signaldetect" value="0" />
-- Retrieval info: 	<generic name="enable_port_rx_std_prbs_status" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="125.0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_clk_network" value="x1" />
-- Retrieval info: </instance>
-- IPFS_FILES : GXB_RX.vho
-- RELATED_FILES: GXB_RX.vhd, altera_xcvr_functions.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_native_av_functions_h.sv, altera_xcvr_native_av.sv, altera_xcvr_data_adapter_av.sv
